--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package constants is

    constant Char_Space : STD_LOGIC_VECTOR(127 downto 0) := (others => '0');
	 constant Char_0 : STD_LOGIC_VECTOR(127 downto 0) :=
	"00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00011100" & 
    "00100010" & 
    "01000101" & 
    "01001001" & 
    "01010001" & 
    "01100001" & 
    "00100010" & 
    "00011100" & 
    "00000000";
	 constant Char_1 : STD_LOGIC_VECTOR(127 downto 0) :=
	 "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00011000" & 
    "00111000" & 
    "01101000" & 
    "00001000" & 
	 "00001000" &
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "01111111" & 
    "00000000";
	 constant Char_2 : STD_LOGIC_VECTOR(127 downto 0) :=
	 "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" &  
    "01111111" & 
    "00000001" & 
	 "00000001" & 
    "00000001" & 
    "01111111" & 
    "01000000" & 
	 "01000000" &
    "01000000" & 
    "01111111" & 
    "00000000";
	 constant Char_3 : STD_LOGIC_VECTOR(127 downto 0) :=
	"00000000"&
	"00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01111111" & 
    "00000001" & 
	 "00000001" & 
    "00000001" & 
    "01111111" & 
    "00000001" &
	 "00000001" & 	 
    "00000001" & 
    "01111111" & 
    "00000000";
	 constant Char_4 : STD_LOGIC_VECTOR(127 downto 0) :=
	 "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01001000" & 
    "01001000" & 
    "01001000" & 
    "01001000" & 
    "01111111" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
	 "00001000" & 
    "00000000";
	 constant Char_5 : STD_LOGIC_VECTOR(127 downto 0) :=
	 "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01111111" & 
    "01000000" & 
    "01000000" & 
	 "01000000" & 
    "01111111" & 
    "00000001" & 
	 "00000001" & 
    "00000001" & 
    "01111111" & 
    "00000000";
	 constant Char_6 : STD_LOGIC_VECTOR(127 downto 0) :=
	 "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" &  
    "01111111" & 
	 "01000000" & 
    "01000000" & 
    "01000000" & 
    "01111111" & 
    "01000001" & 
    "01000001" & 
	 "01000001" &
    "01111111" & 
    "00000000";
	 constant Char_7 : STD_LOGIC_VECTOR(127 downto 0) :=
	 "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01111111" & 
    "00000001" & 
    "00000001" & 
    "00000001" & 
    "00000001" & 
    "00000001" & 
    "00000001" & 
	 "00000001" & 
    "00000001" & 
    "00000000";
	 constant Char_8 : STD_LOGIC_VECTOR(127 downto 0) :=
	 "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01111111" & 
    "01000001" & 
	 "01000001" & 
    "01000001" & 
    "01111111" & 
    "01000001" & 
	 "01000001" & 
    "01000001" & 
    "01111111" & 
    "00000000";
	 constant Char_9 : STD_LOGIC_VECTOR(127 downto 0) :=
	 "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" &  
    "01111111" & 
	 "01000001" & 
    "01000001" & 
    "01000001" & 
    "01111111" & 
    "00000001" & 
	 "00000001" &
    "00000001" & 
    "01111111" & 
    "00000000";

    constant Char_a : STD_LOGIC_VECTOR(127 downto 0) := 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00111100" & 
    "01000010" & 
    "00000010" & 
    "00011110" & 
    "00100010" & 
    "01000010" & 
    "01000110" & 
    "00111011" & 
    "00000000";
    constant Char_b : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "01000000" & 
    "01000000" & 
    "01000000" & 
    "01000000" & 
    "01000000" & 
    "01011100" & 
    "01100010" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01100010" & 
    "01011100" & 
    "00000000";
    constant Char_c : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00011110" & 
    "00100001" & 
    "01000000" & 
    "01000000" & 
    "01000000" & 
    "01000000" & 
    "00100001" & 
    "00011110" & 
    "00000000";
    constant Char_d : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000001" & 
    "00000001" & 
    "00000001" & 
    "00000001" & 
    "00000001" & 
    "00011101" & 
    "00100011" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "00100011" & 
    "00011101" & 
    "00000000";
    constant Char_e : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00011100" & 
    "00100010" & 
    "01000001" & 
    "01111111" & 
    "01000000" & 
    "01000000" & 
    "00100001" & 
    "00011110" & 
    "00000000";
    constant Char_f : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00001100" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "01111100" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00000000";
    constant Char_g : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00011101" & 
    "00100010" & 
    "00100010" & 
    "00011100" & 
    "00100000" & 
    "00111110" & 
    "01000001" & 
    "01000001" & 
    "00111110";
    constant Char_h : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "01000000" & 
    "01000000" & 
    "01000000" & 
    "01000000" & 
    "01000000" & 
    "01011100" & 
    "01100010" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "00000000";
    constant Char_i : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00001000" & 
    "00001000" & 
    "00000000" & 
    "00000000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00000000";
    constant Char_j : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00001000" & 
    "00001000" & 
    "00000000" & 
    "00000000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00110000";
    constant Char_k : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "01000000" & 
    "01000000" & 
    "01000000" & 
    "01000000" & 
    "01000000" & 
    "01000010" & 
    "01000100" & 
    "01001000" & 
    "01010000" & 
    "01101000" & 
    "01000100" & 
    "01000010" & 
    "01000001" & 
    "00000000";
    constant Char_l : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00001000" & 
    "00000000";
    constant Char_m : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01010110" & 
    "01101001" & 
    "01001001" & 
    "01001001" & 
    "01001001" & 
    "01001001" & 
    "01001001" & 
    "01001001" & 
    "00000000";
    constant Char_n : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01011100" & 
    "01100010" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "00000000";
    constant Char_o : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00011100" & 
    "00100010" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "00100010" & 
    "00011100" & 
    "00000000";
    constant Char_p : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01011100" & 
    "01100010" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01100010" & 
    "01011100" & 
    "01000000" & 
    "01000000";
    constant Char_q : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00011101" & 
    "00100011" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "00100011" & 
    "00011101" & 
    "00000001" & 
    "00000001";
    constant Char_r : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00010111" & 
    "00011000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00000000";
    constant Char_s : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00111110" & 
    "01000001" & 
    "01000000" & 
    "00110000" & 
    "00001110" & 
    "00000001" & 
    "01000001" & 
    "00111110" & 
    "00000000";
    constant Char_t : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "01111100" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00010000" & 
    "00001100" & 
    "00000000";
    constant Char_u : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "01000001" & 
    "00100011" & 
    "00011101" & 
    "00000000";
    constant Char_v : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01000001" & 
    "01000001" & 
    "00100010" & 
    "00100010" & 
    "00010100" & 
    "00010100" & 
    "00001000" & 
    "00001000" & 
    "00000000";
    constant Char_w : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01001001" & 
    "01001001" & 
    "01001001" & 
    "01010101" & 
    "01010101" & 
    "00100010" & 
    "00100010" & 
    "00100010" & 
    "00000000";
    constant Char_x : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01000001" & 
    "00100010" & 
    "00010100" & 
    "00001000" & 
    "00001000" & 
    "00010100" & 
    "00100010" & 
    "01000001" & 
    "00000000";
    constant Char_y : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01000001" & 
    "01000001" & 
    "00100010" & 
    "00100010" & 
    "00010100" & 
    "00010100" & 
    "00001000" & 
    "00010000" & 
    "01100000";
    constant Char_z : STD_LOGIC_VECTOR(127 downto 0) :=
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "00000000" & 
    "01111111" & 
    "00000010" & 
    "00000100" & 
    "00001000" & 
    "00010000" & 
    "00100000" & 
    "01000000" & 
    "01111111" & 
    "00000000";

end constants;